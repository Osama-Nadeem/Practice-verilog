module xor(
    a,b,c
)
    input wire a,b;
    output wire c;

    assign c = a ^ b;
endmodule